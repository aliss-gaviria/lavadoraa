library verilog;
use verilog.vl_types.all;
entity lavadora_vlg_vec_tst is
end lavadora_vlg_vec_tst;
